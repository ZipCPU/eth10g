// Goal is to convert from one width to another
//
// Challenges are twofold:
//	1. AXI-Network signaling
//	2. Shift register (not much of a challenge)
//	3. Formal properties
//
// Question: How would you verify this?
// Answer:
//	1. Pick two bytes (like a FIFO). Let them be arbitrary and adjacent.
//		Also, pick their location in the input stream.
//	2. Assume those two bytes arrive on an incoming packet, one after the
//		other.
//	3. *Prove* those same two bytes leave in an outgoing packet, one after
//		the other.
//		Also, *prove* those same two bytes occupy the same locations
//		(byte-wise) in the output stream.
//	4. Assume !S_AXIN_ABORT, *PROVE* !M_AXIN_ABORT
//
`default_nettype none

module	axinwidth #(
        parameter	IW = 64,    // Incoming data path width
        parameter	OW = 32	    // Outgoing data path width
        // Reminder: come back and add these parameters in later
        // parameter [0:0] OPT_LITTLE_ENDIAN
        // parameter [0:0] OPT_LOWPOWER
    ) (
        // {{{
        input	wire					ACLK, ARESETN,
        // S_AXIN_*
        input	wire					S_AXIN_VALID,
        output	wire					S_AXIN_READY,
        input	wire	[IW-1:0]		S_AXIN_DATA,
        input	wire [$clog2(IW/8):0]	S_AXIN_BYTES,
        input	wire					S_AXIN_LAST,
        input	wire					S_AXIN_ABORT,
        // M_AXIN_*
        output	reg		    			M_AXIN_VALID,
        input	wire					M_AXIN_READY,
        output	wire 	[OW-1:0]		M_AXIN_DATA,
        output	reg [$clog2(OW/8):0]	M_AXIN_BYTES,
        output	reg 					M_AXIN_LAST,
        output  reg                     M_AXIN_ABORT
        // }}}
    );

`ifdef FORMAL
    // Pick two arbitrary values
    (* anyconst *) reg	[7:0]	fc_first, fc_next;
    wire	[7:0]	fm_first, fm_next;
    // Pick an arbitrary position
    (* anyconst *) reg	[$clog2(MAX_LENGTH):0]	fc_posn;
    wire	[$clog2(MAX_LENGTH):0]	fc_nxtposn;
`endif

    generate if (IW == OW)
    begin : EQUAL
        // {{{
        assign	S_AXIN_READY = M_AXIN_READY;
        assign	M_AXIN_DATA  = S_AXIN_DATA;
        always @(posedge ACLK) begin
            if (!ARESETN)
            begin
                M_AXIN_VALID <= 0;
                M_AXIN_LAST  <= 0;
                M_AXIN_BYTES <= 0;
                M_AXIN_ABORT <= 0;
            end
            else begin
                M_AXIN_VALID <= S_AXIN_VALID;
                M_AXIN_LAST  <= S_AXIN_LAST;
                M_AXIN_BYTES <= S_AXIN_BYTES;
                M_AXIN_ABORT <= S_AXIN_ABORT;
            end
        end
        // }}}
    end else if (IW < OW)
    // PASSED for ALL
    begin : IW_SMALLER
        // {{{
        // Try IW = 8, OW = 32		(You need this for verification)
        // Also try IW = 32, OW = 64	(I need this for project)
        // Also try IW = 64, OW = 512	(I need this for project)
        integer i;
        localparam SHIFT = IW;
        localparam WIDE_COUNT = (OW/IW);

        reg [OW-1:0] data_concat;
        reg [$clog2(WIDE_COUNT)-1:0] wide_counter;
        reg mid_packet;

        initial mid_packet = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                mid_packet <= 0;
            else if (S_AXIN_ABORT && !S_AXIN_VALID)
                mid_packet <= 0;
            else if (S_AXIN_VALID && S_AXIN_READY)
                mid_packet <= !S_AXIN_LAST && !S_AXIN_ABORT;
        end

        // M_AXIN_ABORT
        initial M_AXIN_ABORT = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                M_AXIN_ABORT <= 0;
            else if (M_AXIN_VALID && !M_AXIN_READY && (M_AXIN_ABORT || (S_AXIN_ABORT && mid_packet)))
                M_AXIN_ABORT <= 1;
            else if (S_AXIN_ABORT && mid_packet)
                M_AXIN_ABORT <= 1;
            else if (!M_AXIN_VALID || M_AXIN_READY)
                M_AXIN_ABORT <= 0;
        end

        // M_AXIN_DATA, S_AXIN_READY
        assign S_AXIN_READY = !M_AXIN_VALID || M_AXIN_READY || S_AXIN_ABORT;
        assign M_AXIN_DATA  = data_concat;

        // M_AXIN_VALID
        initial M_AXIN_VALID = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                M_AXIN_VALID <= 0;
            else begin
                if ((S_AXIN_VALID && S_AXIN_READY) && (wide_counter == WIDE_COUNT-1 || S_AXIN_LAST) && !S_AXIN_ABORT)
                    M_AXIN_VALID <= 1;
                else if (M_AXIN_READY)
                    M_AXIN_VALID <= 0;
            end
        end

        // M_AXIN_BYTES, M_AXIN_LAST, wide_counter, data_concat
        initial M_AXIN_BYTES = 0;
        initial M_AXIN_LAST  = 0;
        initial wide_counter = 0;
        initial data_concat  = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
            begin
                M_AXIN_BYTES <= 0;
                M_AXIN_LAST  <= 0;
                wide_counter <= 0;
                data_concat  <= 0;
            end
            else begin
                if (M_AXIN_VALID && M_AXIN_READY)
                    data_concat <= 0;

                if (S_AXIN_VALID && S_AXIN_READY && !S_AXIN_ABORT)
                begin
                    M_AXIN_LAST <= S_AXIN_LAST;

                    // *_VALID and *_READY can be set at the same time
                    if (M_AXIN_VALID && M_AXIN_READY)
                        M_AXIN_BYTES <= S_AXIN_BYTES;
                    else
                        M_AXIN_BYTES <= M_AXIN_BYTES + S_AXIN_BYTES;

                    for(i=0; i < OW/IW; i=i+1) begin
                        if (wide_counter == i)
                            data_concat[i*IW +: IW] <= S_AXIN_DATA;
                    end

                    if (!S_AXIN_LAST)
                        wide_counter <= wide_counter + 1;
                    else
                        wide_counter <= 0;
                end
                else if ((M_AXIN_VALID && M_AXIN_READY) || (!M_AXIN_VALID && (M_AXIN_ABORT || S_AXIN_ABORT)))
                begin
                    M_AXIN_BYTES <= 0;
                    M_AXIN_LAST  <= 0;
                    wide_counter <= 0;
                    data_concat  <= 0;
                end
            end
        end
        // }}}

////////////////////////////////////////////////////////////////
//
// Formal properties
// {{{
////////////////////////////////////////////////////////////////
`ifdef	FORMAL

    // always @(*) begin
    //     cover(f_m_stream_word == 3);
    // end

    always @(*) begin
        if (ARESETN)
        begin
            if (M_AXIN_VALID && M_AXIN_LAST)
                assert(f_s_stream_word == 0);
            assert(f_m_stream_word < (MAX_LENGTH / (OW/IW)));
            assert(mid_packet == (f_s_stream_word != 0));
            if (!M_AXIN_LAST && !M_AXIN_ABORT)
            begin
                assert(f_m_stream_word <= f_s_stream_word);
                assert(f_s_stream_word == ((f_m_stream_word + (M_AXIN_VALID ? 1:0)) * WIDE_COUNT) + wide_counter);
            end
            assert(!M_AXIN_LAST || M_AXIN_VALID); // ?
            assert(M_AXIN_BYTES <= OW/8);
            if (M_AXIN_BYTES == OW/8)
                assert(M_AXIN_VALID);
            if (!M_AXIN_LAST && !M_AXIN_VALID)
                assert(wide_counter * IW/8 == M_AXIN_BYTES);
            if (M_AXIN_VALID)
                assert(wide_counter == 0);
            assert(data_concat == M_AXIN_DATA);
        end
    end

    assign fm_first = M_AXIN_DATA >> (8*fc_posn[$clog2(OW/8)-1:0]);
    assign fm_next  = M_AXIN_DATA >> (8*fc_nxtposn[$clog2(OW/8)-1:0]);

`endif
// }}}
    end else begin : IW_GREATER // TESTING
        // Try IW=64, OW=32		(I need this for the project)
        // {{{
        integer i;
        localparam PARSE_COUNT = (IW/OW);

        reg shift_en;
        reg [IW-OW-1:0] data_parse;
        reg [$clog2(OW/8):0] remaining_bytes;
        reg remaining_last;
        reg mid_packet;
        reg sready;
        reg [OW-1:0] mdata;

        initial mid_packet = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                mid_packet <= 0;
            else if (S_AXIN_ABORT && !S_AXIN_VALID)
                mid_packet <= 0;
            else if (S_AXIN_VALID && S_AXIN_READY)
                mid_packet <= !S_AXIN_LAST && !S_AXIN_ABORT;
        end

        // M_AXIN_ABORT
        initial M_AXIN_ABORT = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                M_AXIN_ABORT <= 0;
            else if (M_AXIN_VALID && !M_AXIN_READY && (M_AXIN_ABORT || (S_AXIN_ABORT && mid_packet)))
                M_AXIN_ABORT <= 1;
            else if (S_AXIN_ABORT && mid_packet)
                M_AXIN_ABORT <= 1;
            else if (!M_AXIN_VALID || M_AXIN_READY)
                M_AXIN_ABORT <= 0;
        end

        // S_AXIN_READY
        // We shouldn't get the data unless we convey all the incoming data from slave (check!)
        // Don't register s_ready !!!
        // TODO: Add abort here
        assign S_AXIN_READY = !M_AXIN_VALID || (M_AXIN_READY && remaining_bytes == 0);

        // Which word (32-bit) should we send first ?
        // Little endian => sends 0 first
        always @(posedge ACLK) begin
            if (!ARESETN)
                mdata <= 0;
            else if (S_AXIN_VALID && S_AXIN_READY && !S_AXIN_ABORT)
                mdata <= S_AXIN_DATA[0 +: OW];
            else if (M_AXIN_VALID && M_AXIN_READY && !M_AXIN_ABORT)
                mdata <= data_parse[0 +: OW];
        end
        assign M_AXIN_DATA  = mdata;

        // M_AXIN_VALID
        initial M_AXIN_VALID = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
                M_AXIN_VALID <= 0;
            else begin
                if (S_AXIN_VALID && S_AXIN_READY && !S_AXIN_ABORT)
                    M_AXIN_VALID <= 1;
                else if (M_AXIN_READY && (remaining_bytes == 0 || M_AXIN_LAST))
                    M_AXIN_VALID <= 0;
            end
        end

        // M_AXIN_BYTES, M_AXIN_LAST, data_parse
        initial shift_en = 0;
        initial remaining_last = 0;
        initial remaining_bytes = 0;
        initial M_AXIN_BYTES = 0;
        initial M_AXIN_LAST  = 0;
        initial data_parse   = 0;
        always @(posedge ACLK) begin
            if (!ARESETN)
            begin
                shift_en        <= 0;
                remaining_last  <= 0;
                remaining_bytes <= 0;
                M_AXIN_BYTES    <= 0;
                M_AXIN_LAST     <= 0;
                data_parse      <= 0;
            end
            else begin
                if (S_AXIN_VALID && S_AXIN_READY && !S_AXIN_ABORT)
                begin
                    shift_en        <= 0;
                    remaining_bytes <= (S_AXIN_BYTES > OW/8) ? (S_AXIN_BYTES - OW/8) : 0;
                    M_AXIN_BYTES    <= (S_AXIN_BYTES > OW/8) ? (OW/8) : S_AXIN_BYTES[$clog2(OW/8):0];
                    M_AXIN_LAST     <= S_AXIN_LAST && (S_AXIN_BYTES <= OW/8);
                    remaining_last  <= (S_AXIN_LAST && S_AXIN_BYTES > OW/8);
                    data_parse      <= S_AXIN_DATA[IW-1 : OW];
                end
                else if (M_AXIN_VALID && M_AXIN_READY)
                begin
                    shift_en        <= 1;
                    remaining_bytes <= (remaining_bytes <= OW/8) ? 0 : (remaining_bytes - OW/8);
                    M_AXIN_BYTES    <= (remaining_bytes > OW/8) ? OW/8 : remaining_bytes;
                    M_AXIN_LAST     <= (remaining_bytes > OW/8) ? 0 : remaining_last;
                    remaining_last  <= (remaining_bytes <= OW/8) ? 0 : remaining_last;
                    // remaining_last  <= (remaining_bytes <= OW/8) ? 0 : remaining_last;
                    data_parse      <= (shift_en) ? data_parse >> OW : data_parse;
                end
                // else if ((M_AXIN_VALID && M_AXIN_READY) || (!M_AXIN_VALID && (M_AXIN_ABORT || S_AXIN_ABORT)))
                // begin
                //     M_AXIN_BYTES <= 0;
                //     M_AXIN_LAST  <= 0;
                //     data_parse   <= 0;
                // end
            end
        end
        // }}}

////////////////////////////////////////////////////////////////
//
// Formal properties
// {{{
////////////////////////////////////////////////////////////////
`ifdef	FORMAL

    // This one is a challenge to get right, but it is a
    // necessary assertion
    // always @(*)
    //     assert(f_m_stream_word == f_s_stream_word
    //         + (M_AXIN_VALID || (shift_register_valid)));

    always @(*) begin
        cover(f_s_stream_word == 5);
    end

    always @(*) begin
        if (ARESETN)
        begin
            if (M_AXIN_VALID && M_AXIN_LAST)
                assert(f_s_stream_word == 0);
            assert(f_m_stream_word < (MAX_LENGTH * (IW/OW)));
            assert(mid_packet == (f_s_stream_word != 0));
            if (!mid_packet)
                assert(f_s_stream_word == 0);
            if (!mid_packet && !remaining_last && !M_AXIN_LAST)
                assert(f_m_stream_word == 0);
            assert(f_s_stream_word <= f_m_stream_word + 1); // +1 is for first word of slave
            if (mid_packet && remaining_bytes == 0)
                assert((f_s_stream_word * IW/OW) == (f_m_stream_word + (M_AXIN_VALID ? 1:0)));
            assert(M_AXIN_BYTES <= OW/8);
            if (M_AXIN_BYTES == OW/8)
                assert(M_AXIN_VALID);
            if (remaining_bytes > 0)
                assert(!S_AXIN_READY);
            if (mid_packet)
                assert(remaining_last == 0);
        end
    end

    assign fm_first = M_AXIN_DATA >> (8*fc_posn[$clog2(OW/8)-1:0]);
    assign fm_next  = M_AXIN_DATA >> (8*fc_nxtposn[$clog2(OW/8)-1:0]);
`endif
        // }}}
    // }}}
    end endgenerate

////////////////////////////////////////////////////////////////////////////////
//
// Formal properties
// {{{
////////////////////////////////////////////////////////////////////////////////
`ifdef	FORMAL
    localparam MIN_LENGTH = 64*8/IW;
    localparam MAX_LENGTH = 1024;
    localparam LGMX = (MAX_LENGTH > 0) ? $clog2(MAX_LENGTH+1):1;

    // Let the solver pick whether or not we allow aborts
    (* anyconst *) reg	fc_allow_aborts;
    // Pick two arbitrary values
    // (* anyconst *) reg	[IW-1:0]	fc_first, fc_next;
    // wire	[IW-1:0]	fm_first, fm_next;
    // Pick an arbitrary position
    // (* anyconst *) reg	[$clog2(MAX_LENGTH):0]	fc_posn;
    // wire	[$clog2(MAX_LENGTH):0]	fc_nxtposn;

    reg	[LGMX-1:0] f_s_stream_word, f_m_stream_word;
    reg	[12-1:0]   f_s_packets_rcvd, f_m_packets_rcvd;

    reg	f_past_valid;
    initial	f_past_valid = 0;
    always @(posedge ACLK)
        f_past_valid = 1;

    always @(posedge ACLK)
        if (!f_past_valid)
            assume(!ARESETN);

    // fc_nxtposn
    assign	fc_nxtposn = fc_posn + 1;
    always @(*)
    begin
        assume(fc_nxtposn != 0);
        if (S_AXIN_LAST)
            assume(fc_nxtposn < f_s_stream_word);
    end

    ////////////////////////////////////////////////////////////////////////
    //
    // Slave stream properties
    // {{{
    ////////////////////////////////////////////////////////////////////////
    // assume properties of the inputs

    // faxin_slave
    // {{{
    faxin_slave #(
        .DATA_WIDTH(IW),
        .MIN_LENGTH(MIN_LENGTH),
        .MAX_LENGTH(MAX_LENGTH)
    ) fslave (
        .S_AXI_ACLK(ACLK), .S_AXI_ARESETN(ARESETN),
        .S_AXIN_VALID(S_AXIN_VALID),
        .S_AXIN_READY(S_AXIN_READY),
        .S_AXIN_DATA(S_AXIN_DATA),
        .S_AXIN_LAST(S_AXIN_LAST),
        .S_AXIN_ABORT(S_AXIN_ABORT),
        .f_stream_word(f_s_stream_word),
        .f_packets_rcvd(f_s_packets_rcvd)
    );
    // }}}

    // S_AXIN_BYTES
    // {{{
    always @(*) begin
        if (ARESETN && S_AXIN_VALID)
        begin
            assume(S_AXIN_BYTES > 0);
            assume(S_AXIN_BYTES <= IW/8);
            if (!S_AXIN_LAST)
                assume(S_AXIN_BYTES == (IW/8));
        end
    end
    // }}}

    // MIN_LENGTH & S_AXIN_LAST
    // {{{
    always @(*) begin
        if (f_s_stream_word < MIN_LENGTH)
            assume(!S_AXIN_LAST);
    end
    // }}}

    // S_AXIN_ABORT
    // always @(*)
    // if (ARESETN && !fc_allow_aborts)
    //     assume(!S_AXIN_ABORT);

    always @(*)
    if (ARESETN && S_AXIN_VALID && f_s_stream_word == fc_posn[$clog2(MAX_LENGTH):$clog2(IW/8)])
    begin
        // Assume the first data
        if (IW == 8)
            assume(S_AXIN_DATA == fc_first);
        else
            assume(S_AXIN_DATA[fc_posn[$clog2(IW/8)-1:0]*8 +: 8] == fc_first);
    end

    always @(*)
    if (ARESETN && S_AXIN_VALID && f_s_stream_word == fc_nxtposn[$clog2(MAX_LENGTH):$clog2(IW/8)])
    begin
        // Assume the next data
        if (IW == 8)
            assume(S_AXIN_DATA == fc_next);
        else
            assume(S_AXIN_DATA[fc_nxtposn[$clog2(IW/8)-1:0]*8 +: 8] == fc_next);
    end
    // }}}

    ////////////////////////////////////////////////////////////////////////
    //
    // Master stream properties
    // {{{
    ////////////////////////////////////////////////////////////////////////
    // assert properties of the outputs

    // faxin_master
    faxin_master #(
        .DATA_WIDTH(OW),
        .MIN_LENGTH(MIN_LENGTH*(IW/OW)),
        .MAX_LENGTH(MAX_LENGTH*(IW/OW))
    ) fmaster (
        .S_AXI_ACLK(ACLK), .S_AXI_ARESETN(ARESETN),
        .S_AXIN_VALID(M_AXIN_VALID),
        .S_AXIN_READY(M_AXIN_READY),
        .S_AXIN_DATA(M_AXIN_DATA),
        .S_AXIN_LAST(M_AXIN_LAST),
        .S_AXIN_ABORT(M_AXIN_ABORT),
        .f_stream_word(f_m_stream_word),
        .f_packets_rcvd(f_m_packets_rcvd)
    );

    // M_AXIN_ABORT
    // always @(*)
    // if (ARESETN && !fc_allow_aborts)
    //     assert(!M_AXIN_ABORT);

    always @(*)
    if (ARESETN && M_AXIN_ABORT)
        assert(f_s_stream_word == 0);

    always @(*)
    if (ARESETN && !M_AXIN_ABORT && (f_s_stream_word > (fc_posn[$clog2(MAX_LENGTH):$clog2(IW/8)]) || M_AXIN_LAST)
        && f_m_stream_word == fc_posn[$clog2(MAX_LENGTH):$clog2(OW/8)])
    begin
        // Assert the first data
        assert(fm_first == fc_first);
    end

    always @(*)
    if (ARESETN && !M_AXIN_ABORT && (f_s_stream_word > (fc_nxtposn[$clog2(MAX_LENGTH):$clog2(IW/8)]) || M_AXIN_LAST)
        && f_m_stream_word == fc_nxtposn[$clog2(MAX_LENGTH):$clog2(OW/8)])
    begin
        // Assert the next data
        assert(fm_next == fc_next);
    end

    // M_AXIN_BYTES
    // {{{
    always @(*)
    if (M_AXIN_VALID)
    begin
        assert(M_AXIN_BYTES > 0);
        assert(M_AXIN_BYTES <= OW/8);
        if (!M_AXIN_LAST)
            assert(M_AXIN_BYTES == OW/8);
    end
    // }}}

    // }}}
    ////////////////////////////////////////////////////////////////////////
    //
    // Low power rules (if we wish to use them
    // {{{
    ////////////////////////////////////////////////////////////////////////

    /*
    // Power is used every time a register toggles
    // So, if OPT_LOWPOWER is set -- we keep registers from toggling
    //	(by pinning them to zero)
    always @(*)
    if (OPT_LOWPOWER && !M_AXIN_VALID)
    begin
        // Can't assert these first two, since you are building
        // in M_AXIN_DATA while !M_AXIN_VALID, so we won't assert
        // these at all.
        //
        // assert(M_AXIN_DATA  == 0);
        // assert(M_AXIN_BYTES == 0);
        //

        if (WIDE_COUNT == 0)
            assert(M_AXIN_DATA == 0);

        assert(M_AXIN_LAST  == 0);
    end

    always @(*)
    if (OPT_LOWPOWER && M_AXIN_VALID)
    begin
        for(i=0; i<OW/8; i=i+1)
        if (i >= M_AXIN_BYTES)
            assert(M_AXIN_DATA[8*i +: 8] == 0);
    end
    */
    // }}}
    ////////////////////////////////////////////////////////////////////////
    //
    // "Careless" assumptions
    // {{{
    ////////////////////////////////////////////////////////////////////////
    //
    //

    // Just to get us started, and give us some confidence that this is
    // working
    always @(*)
        assume(!S_AXIN_ABORT);

    // }}}
`endif
// }}}
endmodule
