../../wbsata/rtl/sata_primitives.vh